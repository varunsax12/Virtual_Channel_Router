
`ifndef VR_define
`define VR_define

`define MATRIX_ARBITER        1
`define ROUND_ROBIN_ARBITER   2

`define ARBITER_TYPE          2

`endif