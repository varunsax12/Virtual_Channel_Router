
`ifndef VR_define
`define VR_define

`define MATRIX_ARBITER        1
`define ROUND_ROBIN_ARBITER   2

`define SEPARABLE_ALLOCATOR   1
`define WAVEFRONT_ALLOCATOR   2

`define ARBITER_TYPE          1

`define ALLOCATOR_TYPE        1

`endif
